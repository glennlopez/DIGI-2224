-- set library
library ieee;

-- set entity as filename

-- set architechture
	-- set select statement
