library verilog;
use verilog.vl_types.all;
entity truth_table_1_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end truth_table_1_vlg_check_tst;
