library ieee;use ieee.std_logic_1164.all;use ieee.std_logic_arith.all;entity full_adder_tb isend full_adder_tb;architecture test_bench of full_adder_tb is	component full_adder		port		(			a, b, c_in : in std_logic;			c_out, sum : out std_logic		);	end component;	signal operands : std_logic_vector(2 downto 0);signal result : std_logic_vector(1 downto 0);beginfull_add: full_adder port map( a => operands(2),b => operands(1),c_in => operands(0),c_out => result(1),sum => result(0));stim_proc: processbeginfor j in 0 to 7 loopoperands <= CONV_STD_LOGIC_VECTOR(j,3);wait for 100 ns;end loop;wait;end process;end test_bench;