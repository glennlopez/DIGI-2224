library verilog;
use verilog.vl_types.all;
entity truth_table_1_vlg_vec_tst is
end truth_table_1_vlg_vec_tst;
