-- set library

-- set entity as filename

-- set architechture
	-- set select statement
