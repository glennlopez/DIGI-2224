-- full_adder_tb.vhd-- test bench for full_adder.vhd-- simulation criteria:-- 2-bit output = sum of three 1-bit inputs-- Test by applying a binary count on the inputslibrary ieee;use ieee.std_logic_1164.all;use ieee.std_logic_arith.all;entity full_adder_tb is-- test bench entity has no external portsend full_adder_tb;architecture test_bench of full_adder_tb iscomponent full_adderport(a, b, c_in : in std_logic;c_out, sum : out std_logic);end component;signal operands : std_logic_vector(2 downto 0);signal result : std_logic_vector(1 downto 0);begin-- instantiate full adder with test signalsfull_add: full_adder port map( a => operands(2),b => operands(1),c_in => operands(0),c_out => result(1),sum => result(0));-- stimulus process (generates simulation input waveforms)stim_proc: processbegin-- Count from 0 to 7for j in 0 to 7 loop-- Convert integer count to 3-bit std_logic_vectoroperands <= CONV_STD_LOGIC_VECTOR(j,3);-- Set time interval for each input statewait for 100 ns;end loop;wait; -- stall here (simulation done)end process;end test_bench;