----------------------------------------------------------------------
--			LAB4: quad2to1.vhd
--
--		Write a VHDL file that defines a multiplexer that switches 
--		two 4-bit inputs, x and y to a 4-bit output, z. Define x, y, 
--		and z as type BIT_VECTOR
----------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

--entity
entity quad2to1 is
  port (
	
  );
end entity;

--architecture

